* draft7
r12 1 2 1.2
r23 2 3 2.3
r1 1 ITerm1 1e-3
r2 2 ITerm2 1e-3
r3 ITerm3 3 1e-3
i1 ITerm1 0 1
i2 ITerm2 0 2
i3 ITerm3 0 3
v1 1 0 1
v2 2 0 2
v3 3 0 3
.op
.backanno
.end
