* draft6

* Resistive network
R0 n00 n01 1.25
R1 n01 n02 1.25
R2 n02 n03 1.25
R3 n10 n11 1.25
R4 n11 n12 1.25
R5 n12 n13 1.25
R6 n20 n21 1.25
R7 n21 n22 1.25
R8 n22 n23 1.25
R9 n30 n31 1.25
R10 n31 n32 1.25
R11 n32 n33 1.25
R12 n00 n10 1.25
R13 n10 n20 1.25
R14 n20 n30 1.25
R15 n01 n11 1.25
R16 n11 n21 1.25
R17 n21 n31 1.25
R18 n02 n12 1.25
R19 n12 n22 1.25
R20 n22 n32 1.25
R21 n03 n13 1.25
R22 n13 n23 1.25
R23 n23 n33 1.25

* Sinks
I0 n00 0 0.3125m
I1 n01 0 0.3125m
I2 n02 0 0.3125m
I3 n03 0 0.3125m
I4 n10 0 0.3125m
I5 n11 0 0.3125m
I6 n12 0 0.3125m
I7 n13 0 0.3125m
I8 n20 0 0.3125m
I9 n21 0 0.3125m
I10 n22 0 0.3125m
I11 n23 0 0.3125m
I12 n30 0 0.3125m
I13 n31 0 0.3125m
I14 n32 0 0.3125m
I15 n33 0 0.3125m

* Sources
V0 n00 0 1.8
V1 n01 0 1.8
V2 n02 0 1.8
V3 n03 0 1.8
V4 n10 0 1.8
V5 n11 0 1.8
V6 n12 0 1.8
V7 n13 0 1.8
V8 n20 0 1.8
V9 n21 0 1.8
V10 n22 0 1.8
V11 n23 0 1.8
V12 n30 0 1.8
V13 n31 0 1.8
V14 n32 0 1.8
V15 n33 0 1.8

*Footer
.OPTION NUMDGT=6
.OP
.SAVE TYPE=IC FILE=compare.ic
.END
