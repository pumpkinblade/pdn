* draft7
r12 1 2 0.5
r23 2 3 0.25
i1 1 0 1
i2 2 0 2
i3 3 0 3
r1 1 x1 0.1
r2 2 x2 0.1
r3 3 x3 0.1
v1 x1 0 1
v2 x2 0 2
v3 x3 0 3
.op
.backanno
.end
